p(X) :- q(X) :0.3.
p(X) :- r(X), p(X) :0.3.
q(1) :1.0.
r(1) :1.0.