p(X,Y) :- edge(X,Y) : 0.5.
p(X,Z) :- p(X,Y), p(Y,Z) : 0.5.
edge(0, 1): 0.5.
edge(1, 0): 0.5.