p(X,Y) :- edge(X,Y) : 0.5.

p(X,Z) :- p(X,Y), p(Y,Z) : 0.5.

edge(0, 1): 0.5.

edge(1, 2): 0.5.

edge(2, 3): 0.5.

edge(3, 4): 0.5.

edge(4, 5): 0.5.

edge(5, 0): 0.5.