p(X,Y) :-e(X,Z), e(Z,Y).
e(0,1).
e(1,2).