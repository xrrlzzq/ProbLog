p(X,Y) :- e(X,Y) :0.5.
p(X,Y) :- e(X,Z), p(Z,Y) :0.5.
e(1,2) :0.5.
e(2,3) :0.5.
e(3,4) :0.5.
e(4,5) :0.5.
e(5,1) :0.5.