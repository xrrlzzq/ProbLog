p(X,Y) :- edge(X,Y) : 0.5.
p(X,Z) :- edge(X,Y), p(Y,Z) : 0.5.
edge(0, 1): 0.5.
edge(1, 2): 0.5.
edge(2, 3): 0.5.
edge(3, 4): 0.5.
edge(4, 5): 0.5.
edge(5, 6): 0.5.
edge(6, 7): 0.5.
edge(7, 8): 0.5.
edge(8, 9): 0.5.
edge(9, 10): 0.5.
edge(10, 11): 0.5.
edge(11, 12): 0.5.
edge(12, 13): 0.5.
edge(13, 14): 0.5.
edge(14, 15): 0.5.
edge(15, 16): 0.5.
edge(16, 17): 0.5.
edge(17, 18): 0.5.
edge(18, 19): 0.5.
edge(19, 20): 0.5.
edge(20, 21): 0.5.
edge(21, 22): 0.5.
edge(22, 23): 0.5.
edge(23, 24): 0.5.
edge(24, 25): 0.5.
edge(25, 26): 0.5.
edge(26, 27): 0.5.
edge(27, 28): 0.5.
edge(28, 29): 0.5.
edge(29, 30): 0.5.
edge(30, 31): 0.5.
edge(31, 32): 0.5.
edge(32, 33): 0.5.
edge(33, 34): 0.5.
edge(34, 35): 0.5.
edge(35, 36): 0.5.
edge(36, 37): 0.5.
edge(37, 38): 0.5.
edge(38, 39): 0.5.
edge(39, 40): 0.5.
edge(40, 41): 0.5.
edge(41, 42): 0.5.
edge(42, 43): 0.5.
edge(43, 44): 0.5.
edge(44, 45): 0.5.
edge(45, 46): 0.5.
edge(46, 47): 0.5.
edge(47, 48): 0.5.
edge(48, 49): 0.5.
edge(49, 50): 0.5.