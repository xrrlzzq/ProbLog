p(X,Y) :- e(X,Y) :0.8.
p(X,Z) :- e(X,Z), e(Z,Y) :0.6.
e(2,1) :0.7.
e(2,4) :0.3.
e(1,4) :0.1.
e(3,2) :0.5.