p(X,Y):-e(X,Y).
p(X,Y):-p(X,Z),p(Z,Y).
e(1,2).
e(2,3).
e(3,1).
e('a B',1).