p(X,Y) :- e(X,Y) :0.8.
p(X,Z) :- e(X,Z), p(X,Y) :0.6.
e(0,1) :0.5.
e(0,2) :0.7.
e(1,3) :0.3.