p(X,Y) :- p(X,Y), q(Y,Z) : 0.3.
p(0,1): 0.5.
q(1,2): 0.3.